library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity keypad_logic is
--  Port ( );
end keypad_logic;

architecture Behavioral of keypad_logic is

begin


end Behavioral;
