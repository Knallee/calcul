library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity edge_det is
--  Port ( );
end edge_det;

architecture Behavioral of edge_det is

begin


end Behavioral;
