library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity keypad_top is
--  Port ( );
end keypad_top;

architecture Behavioral of keypad_top is

begin


end Behavioral;
