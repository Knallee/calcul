library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity debouncer is
--  Port ( );
end debouncer;

architecture Behavioral of debouncer is

begin


end Behavioral;
